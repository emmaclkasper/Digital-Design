`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: Courtney Trust and Emma Kasper
// 
// Create Date:    12:46:07 10/17/2019 
// Design Name: 
// Module Name:    Binary2BCD_tb 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module Binary2BCD_tb();

	reg [3:0]Cnt_s;
	wire [3:0]Tens_s, Ones_s;
	
	Binary2BCD ComptoTest(Cnt_s, Tens_s, Ones_s);
	
	//Vector Procedure
	initial begin
		#10 Cnt_s <= 4'b0000;
		#10 Cnt_s <= 4'b0001;
		#10 Cnt_s <= 4'b0010;
		#10 Cnt_s <= 4'b0011;
		#10 Cnt_s <= 4'b0100;
		#10 Cnt_s <= 4'b0101;
		#10 Cnt_s <= 4'b0110;
		#10 Cnt_s <= 4'b0111;
		#10 Cnt_s <= 4'b1000;
		#10 Cnt_s <= 4'b1001;
		#10 Cnt_s <= 4'b1010;
		#10 Cnt_s <= 4'b1011;
		#10 Cnt_s <= 4'b1100;
		#10 Cnt_s <= 4'b1101;
		#10 Cnt_s <= 4'b1110;
		#10 Cnt_s <= 4'b1111;
	
	end

endmodule
